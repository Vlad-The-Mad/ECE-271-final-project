module RAM (input logic [15:0] read_address,
            input logic [15:0] write_address,
            input logic [15:0] write_value,
            output logic [15:0] word);

endmodule
